
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;

entity InstructionMemory is 
    generic (
        PC_WIDTH  : integer := 32;  -- instruction width 
        MEM_DEPTH : integer := 128   -- instruction depth 
    );
    port (
        i_address     : in std_ulogic_vector(PC_WIDTH-1 downto 0);
        o_instruction : out std_ulogic_vector(PC_WIDTH-1 downto 0)
    );
end entity InstructionMemory;

architecture RTL of InstructionMemory is 
    signal index : integer := 0;
    type memory_array is array (0 to MEM_DEPTH-1) of std_ulogic_vector(PC_WIDTH-1 downto 0);

    constant instruction_array : memory_array := (
        0   => x"00000013",  
        1   => x"00000093",  
        2   => x"002081B3",  
        3   => x"403181B3",  
        4   => x"00209233",  
        5   => x"0020A2B3",  
        6   => x"0020B333",  
        7   => x"0020C3B3",  
        8   => x"0020D433",  
        9   => x"4020D433",
        10  => x"0020E4B3", 
        11  => x"0020F533", 
        12  => x"00210113",
        13  => x"00310193", 
        14  => x"00418213", 
        15  => x"00520293", 
        16  => x"00628313", 
        17  => x"00730393", 
        18  => x"00838413", 
        19  => x"40840493", 
        20  => x"00948513", 
        21  => x"00A50593", 
        22  => x"00058663", 
        23  => x"00160663", 
        24  => x"00268663", 
        25  => x"00370663", 
        26  => x"00478663", 
        27  => x"00580663", 
        28  => x"0000006F", 
        29  => x"000080E7", 
        30  => x"00002003", 
        31  => x"00113003", 
        32  => x"00214003", 
        33  => x"00315003", 
        34  => x"00416003", 
        35  => x"00512023", 
        36  => x"00613023", 
        37  => x"00714023", 
        38  => x"020000F3", 
        39  => x"020080F3", 
        40  => x"0200C0F3", 
        41  => x"0201C0F3", 
        42  => x"020140F3", 
        43  => x"0202C0F3", 
        44  => x"020340F3", 
        45  => x"020440F3", 
        46  => x"0204C0F3", 
        47  => x"020540F3", 
        48  => x"0205C0F3", 
        49  => x"000200B3", 
        50  => x"000240B3", 
        51  => x"000280B3", 
        52  => x"0002C0B3", 
        53  => x"000300B3", 
        54  => x"000340B3", 
        55  => x"000380B3", 
        56  => x"0003C0B3", 
        57  => x"00000073", 
        58  => x"00100073", 
        59  => x"0000100F", 
        60  => x"0000100F",
        61  => x"00000013",  
        62  => x"00000093",  
        63  => x"002081B3",  
        64  => x"00209233",  
        65  => x"0020A2B3",  
        66  => x"0020B333",  
        67  => x"0020C3B3",  
        68  => x"0020D433",  
        69  => x"4020D433",
        70  => x"0020E4B3", 
        71  => x"0020F533", 
        72  => x"00210113",
        73  => x"00310193", 
        74  => x"00418213", 
        75  => x"00520293", 
        76  => x"00628313", 
        77  => x"00730393", 
        78  => x"00838413", 
        79  => x"40840493", 
        80  => x"00948513", 
        81  => x"00A50593", 
        82  => x"00058663", 
        83  => x"00160663", 
        84  => x"00268663", 
        85  => x"00370663", 
        86  => x"00478663", 
        87  => x"00580663", 
        88  => x"0000006F", 
        89  => x"000080E7", 
        90  => x"00002003", 
        91  => x"00113003", 
        92  => x"00214003", 
        93  => x"00315003", 
        94  => x"00416003", 
        95  => x"00512023", 
        96  => x"00613023", 
        97  => x"00714023", 
        98  => x"020000F3", 
        99  => x"020080F3", 
        100 => x"0200C0F3", 
        101 => x"0201C0F3", 
        102 => x"020140F3", 
        103 => x"0202C0F3", 
        104 => x"020340F3", 
        105 => x"020440F3", 
        106 => x"0204C0F3", 
        107 => x"020540F3", 
        108 => x"0205C0F3", 
        109 => x"000200B3", 
        110 => x"000240B3", 
        111 => x"000280B3", 
        112 => x"0002C0B3", 
        113 => x"000300B3", 
        114 => x"000340B3", 
        115 => x"000380B3", 
        116 => x"0003C0B3", 
        117 => x"00000073", 
        118 => x"00100073", 
        119 => x"0000100F", 
        120 => x"0000100F",
        121 => x"403181B3",
        122 => x"020140F3", 
        123 => x"0202C0F3", 
        124 => x"020340F3", 
        125 => x"020440F3", 
        126 => x"0204C0F3", 
        127 => x"020540F3",
        others => x"00000000"
    );
    begin 
    process(i_address) is 
        begin 
            index <= to_integer(unsigned(i_address(31 downto 2)));
            if (index < MEM_DEPTH) then 
                o_instruction <= instruction_array(index);
            else 
                o_instruction <= (others => '0'); -- NOP 
            end if;
    end process;
end architecture RTL;


